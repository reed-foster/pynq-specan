../../audio_visualizer_rgb.srcs/sources_1/new/adau1761.sv