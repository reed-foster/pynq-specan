../../audio_visualizer_rgb.srcs/sources_1/new/sample_buffer.sv