../../audio_visualizer_rgb.srcs/sources_1/new/ws2812b.sv