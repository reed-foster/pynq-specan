../../audio_visualizer_rgb.srcs/sources_1/new/axis.sv