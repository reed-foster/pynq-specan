../../audio_visualizer_rgb.srcs/sources_1/new/psd_estimator.sv